module vga_draw(
	input clk,
	input rst,
	input [9:0] x_coord,
	input [9:0] y_coord,
	input video_on,
	input [9:0] start_x,
	input [9:0] start_y,
	input [9:0]end_x,
	input [9:0]end_y,
	input [23:0] bkg_rgb,
	output reg shape_active
	);
	
endmodule